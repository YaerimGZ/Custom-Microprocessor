-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: miche
-- 
-- Create Date:    02/06/2021 00:32:25
-- Project Name:   MEMORIA
-- Module Name:    MEMORIA.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;  -- Para std_logic
use IEEE.numeric_std.all;     -- Para unsigned

entity MEMORIA is
	port(A: IN STD_LOGIC_VECTOR(8 downto 0);
		D: INOUT STD_LOGIC_VECTOR(7 downto 0);
		WR, OE, CS: IN STD_LOGIC);
end MEMORIA;

architecture arq1 of MEMORIA is

	type RAM is array (0 to 511) of std_logic_vector(7 downto 0);
	signal contenido : RAM := (x"84",x"06",x"04",x"08",x"D6",x"F0",x"D9",x"FA",
   			  				   x"29",x"DC",x"F0",x"DB",x"FB",x"9C",x"00",x"00",
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",	
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		

   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",	
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",			

   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",	
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",	

   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",	
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",		
   			  				   x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");

	signal palabra: integer range 0 to 511 := 0;
begin
	process (A, D, WR, OE, CS, contenido, palabra)
		begin
			palabra <= to_integer(unsigned(A(8 downto 0)));
				if OE = '0' and CS = '0' then
					D <= contenido(palabra);
				elsif WR = '0' and CS = '0' then
					contenido(palabra) <= D;
				else
					D <= "ZZZZZZZZ";
				end if;

end process;

end arq1;
