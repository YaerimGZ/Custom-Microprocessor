-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: miche
-- 
-- Create Date:    02/06/2021 00:08:33
-- Project Name:   CONTROL
-- Module Name:    CONTROL.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;  -- Para std_logic
use IEEE.numeric_std.all;     -- Para unsigned

entity CONTROL is
	port(COOP: IN STD_LOGIC_VECTOR(7 downto 0);
		RESET, CLK: IN STD_LOGIC;
		SCONTROL: OUT STD_LOGIC_VECTOR(15 downto 0));
end CONTROL;

architecture arq1 of CONTROL is
	type ROM is array (0 to 1791) of STD_LOGIC_VECTOR(15 downto 0);
	signal CONTENIDO : ROM := ( x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B4", x"00B8", x"00B8",--SUM #,R1
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8",--SUM R1, R1
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8",--SUM R2, R1
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8",--SUM R3, R1
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B2", x"00B8", x"00B8",--SUM #, R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8",--SUM R1, R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8",--SUM R2, R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8",--SUM R3, R2
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B1", x"00B8", x"00B8",--SUM #, R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8",--SUM R1, R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8",--SUM R2, R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8",--SUM R3, R3

								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"14b8", x"0198", x"00B4", x"00B8", x"00B8",--RES # R1
								x"14B8", x"0198", x"0078", x"0078", x"00B4", x"00B8", x"00B8", x"00B8",--RES R1,R1
								x"14B8", x"0198", x"0078", x"0078", x"00B4", x"00B8", x"00B8", x"00B8",--RES R2,R1
								x"14B8", x"0198", x"0078", x"0078", x"00B4", x"00B8", x"00B8", x"00B8",--RES R3,R1
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B2", x"00B8", x"00B8",--RES #,R2
								x"14B8", x"0198", x"0078", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", --RES R1,R2
								x"14B8", x"0198", x"0078", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", --RES R2,R2
								x"14B8", x"0198", x"0078", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", --RES R3, R2
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B1", x"00B8", x"00B8", --RES #, R3
								x"14B8", x"0198", x"0078", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", --RES R1,R3
								x"14B8", x"0198", x"0078", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", --RES R2,R3
								x"14B8", x"0198", x"0078", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", --RES R3, R3

								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B4", x"00B8", x"00B8", --MUL #, R1
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --MUL R1, R1
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --MUL R2, R1
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --MUL R3, R1
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B2", x"00B8", x"00B8", --MUL #, R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --MUL R1, R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --MUL R2, R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --MUL R3, R2
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B1", x"00B8", x"00B8", --MUL #, R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --MUL R1, R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --MUL R2, R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --MUL R3, R3

								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B4", x"00B8", x"00B8", --DIV #, R1
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --DIV R1, R1 
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --DIV R2, R1
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --DIV R3, R1
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B2", x"00B8", x"00B8", --DIV #, R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --DIV R1, R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --DIV R2, R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --DIV R3, R2
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B1", x"00B8", x"00B8", --DIV #, R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --DIV R1, R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --DIV R2, R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --DIV R3, R3

								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B4", x"00B8", x"00B8", --AND #, R1
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --AND R1, R1
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --AND R2, R1
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --AND R3, R1
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B2", x"00B8", x"00B8", --AND #, R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --AND R1, R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --AND R2, R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --AND R3, R2
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B1", x"00B8", x"00B8", --AND #, R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --AND R1, R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --AND R2, R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --AND R3, R3

								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B4", x"00B8", x"00B8", --OR #,R1
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --OR R1,R1 
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --OR R2,R1 
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --OR R3,R1
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B2", x"00B8", x"00B8", --OR #,R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --OR R1,R2 
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --OR R2,R2 
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --OR R3,R2
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B1", x"00B8", x"00B8", --OR #,R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --OR R1,R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --OR R2,R3 
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --OR R3,R3
 
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --NOT R1 
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --NOT R2 
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --NOT R3
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --IZQ R1 
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --IZQ R2 
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --IZQ R3
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --DER R1 
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --DER R2 
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --DER R3
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",

								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B4", x"00B8", x"00B8", --XOR #,R1
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --XOR R1,R1 
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --XOR R2,R1 
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --XOR R3,R1
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B2", x"00B8", x"00B8", --XOR #,R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --XOR R1,R2 
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --XOR R2,R2 
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --XOR R3,R2
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B1", x"00B8", x"00B8", --XOR #,R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --XOR R1,R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --XOR R2,R3 
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --XOR R3,R3 

								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B4", x"00B8", x"00B8", --MOV #,R1
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --MOV R1,R3
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --MOV R2,R3 
								x"14B8", x"0198", x"0078", x"00B4", x"00B8", x"00B8", x"00B8", x"00B8", --MOV R3,R3 
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B2", x"00B8", x"00B8", --MOV #,R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --MOV R1,R2
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --MOV R2,R2 
								x"14B8", x"0198", x"0078", x"00B2", x"00B8", x"00B8", x"00B8", x"00B8", --MOV R3,R2 
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B1", x"00B8", x"00B8", --MOV #,R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --MOV R1,R3
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --MOV R2,R3 
								x"14B8", x"0198", x"0078", x"00B1", x"00B8", x"00B8", x"00B8", x"00B8", --MOV R3,R3

								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --MAY DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --MAY DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --MAY DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --MAY DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --MEN DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --MEN DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --MEN DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --MEN DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --EQU DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --EQU DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --EQU DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --EQU DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --INC DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --INC DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --INC DIR
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0938", x"00B8", x"00B8", --INC DIR

								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",

								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",

								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B0", x"00B8", x"00B8", --COMP R1,X
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B0", x"00B8", x"00B8", --COMP R2,X
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B0", x"00B8", x"00B8", --COMP R3,X
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B0", x"00B8", x"00B8", --COMP R1,R1
								x"14B8", x"0198", x"0078", x"00B0", x"00B8", x"00B8", x"00B8", x"00B8", --COMP R1,R1
								x"14B8", x"0198", x"0078", x"00B0", x"00B8", x"00B8", x"00B8", x"00B8", --COMP R2,R1
								x"14B8", x"0198", x"0078", x"00B0", x"00B8", x"00B8", x"00B8", x"00B8", --COMP R3,R1
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B0", x"00B8", x"00B8", --COMP X,R2
								x"14B8", x"0198", x"0078", x"00B0", x"00B8", x"00B8", x"00B8", x"00B8", --COMP R1,R2
								x"14B8", x"0198", x"0078", x"00B0", x"00B8", x"00B8", x"00B8", x"00B8", --COMP R2,R2
								x"14B8", x"0198", x"0078", x"00B0", x"00B8", x"00B8", x"00B8", x"00B8", --COMP R3,R2
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"00B0", x"00B8", x"00B8", --COMP X,R3
								x"14B8", x"0198", x"0078", x"00B0", x"00B8", x"00B8", x"00B8", x"00B8", --COMP R1,R3
								x"14B8", x"0198", x"0078", x"00B0", x"00B8", x"00B8", x"00B8", x"00B8", --COMP R2,R3
								x"14B8", x"0198", x"0078", x"00B0", x"00B8", x"00B8", x"00B8", x"00B8", --COMP R3,R3

								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8",
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0638", x"019C", x"019C", --MOV X,R1
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0638", x"019C", x"019C", --MOV X,R1
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0638", x"00A0", x"00A0", --MOV R1,X
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0638", x"00A0", x"00A0", --MOV R1,X
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0638", x"019A", x"019A", --MOV X,R2
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0638", x"019A", x"019A", --MOV X,R2
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0638", x"00A0", x"00A0", --MOV R2,X
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0638", x"00A0", x"00A0", --MOV R2,X
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0638", x"0199", x"0199", --MOV X,R3
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0638", x"0199", x"0199", --MOV X,R3
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0638", x"00A0", x"00A0", --MOV R3,X
								x"14B8", x"0198", x"0078", x"14B8", x"0198", x"0638", x"00A0", x"00A0"  --MOV R3,X
			);

	signal PALABRA: integer range 0 to 1791 := 0;
	signal CONTADOR: STD_LOGIC_VECTOR(2 downto 0) := "000";
	signal DIRECCION: STD_LOGIC_VECTOR(10 downto 0);

begin

	process(COOP, RESET, CLK)
		variable TEMPCONT : unsigned(2 downto 0):= "000";

		begin
			if CLK'event and CLK = '1' then
				if RESET = '0' then
						TEMPCONT := "000";
				else
					TEMPCONT := TEMPCONT + 1;
				end if;
			end if;
		CONTADOR <= STD_LOGIC_VECTOR(TEMPCONT);
	end process;

	DIRECCION <= COOP & CONTADOR;
	PALABRA <= TO_INTEGER(UNSIGNED(DIRECCION));
	SCONTROL <= CONTENIDO(PALABRA);


end arq1;
